module vector_dot_prod(
    vec_a_0, vec_a_1, vec_a_2, vec_a_3,
    vec_b_0, vec_b_1, vec_b_2, vec_b_3,
    product_0, product_1, product_2, product_3
    );

